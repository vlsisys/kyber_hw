// ==================================================
//	[ VLSISYS Lab. ]
//	* Author		: Woong Choi (woongchoi@sm.ac.kr)
//	* Filename		: cbd.v
//	* Description	: 
// ==================================================

module cbd
(	
	output reg	[256*4-1:0]		o_coeff,
	input		[64*8-1:0]		i_ibytes,
	input		[1:0]			i_eta
);



endmodule
